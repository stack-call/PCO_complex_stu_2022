library verilog;
use verilog.vl_types.all;
entity cpu is
    port(
        data_in         : in     vl_logic_vector(7 downto 0);
        clk_quick       : in     vl_logic;
        clk_slow        : in     vl_logic;
        clk_delay       : in     vl_logic;
        rst             : in     vl_logic;
        SW_choose       : in     vl_logic;
        A1              : in     vl_logic;
        cpustate        : in     vl_logic_vector(1 downto 0);
        addr            : out    vl_logic_vector(15 downto 0);
        data_out        : out    vl_logic_vector(7 downto 0);
        r0dbus          : out    vl_logic_vector(7 downto 0);
        r1dbus          : out    vl_logic_vector(7 downto 0);
        zout            : out    vl_logic;
        read            : out    vl_logic;
        write           : out    vl_logic;
        arload          : out    vl_logic;
        arinc           : out    vl_logic;
        pcinc           : out    vl_logic;
        pcload          : out    vl_logic;
        drload          : out    vl_logic;
        trload          : out    vl_logic;
        irload          : out    vl_logic;
        r1load          : out    vl_logic;
        r0load          : out    vl_logic;
        xload           : out    vl_logic;
        zload           : out    vl_logic;
        pcbus           : out    vl_logic;
        drhbus          : out    vl_logic;
        drlbus          : out    vl_logic;
        trbus           : out    vl_logic;
        r1bus           : out    vl_logic;
        r0bus           : out    vl_logic;
        membus          : out    vl_logic;
        busmem          : out    vl_logic;
        clr             : out    vl_logic
    );
end cpu;
