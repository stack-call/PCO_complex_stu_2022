library verilog;
use verilog.vl_types.all;
entity light_show is
    port(
        light_clk       : in     vl_logic;
        SW_choose       : in     vl_logic;
        check_in        : in     vl_logic_vector(7 downto 0);
        read            : in     vl_logic;
        write           : in     vl_logic;
        arload          : in     vl_logic;
        arinc           : in     vl_logic;
        pcinc           : in     vl_logic;
        pcload          : in     vl_logic;
        drload          : in     vl_logic;
        trload          : in     vl_logic;
        irload          : in     vl_logic;
        r1load          : in     vl_logic;
        r0load          : in     vl_logic;
        zload           : in     vl_logic;
        pcbus           : in     vl_logic;
        drhbus          : in     vl_logic;
        drlbus          : in     vl_logic;
        trbus           : in     vl_logic;
        r1bus           : in     vl_logic;
        r0bus           : in     vl_logic;
        membus          : in     vl_logic;
        busmem          : in     vl_logic;
        clr             : in     vl_logic;
        State           : in     vl_logic_vector(1 downto 0);
        MAR             : in     vl_logic_vector(7 downto 0);
        r0              : in     vl_logic_vector(7 downto 0);
        r1              : in     vl_logic_vector(7 downto 0);
        Z               : in     vl_logic;
        HEX0            : out    vl_logic_vector(6 downto 0);
        HEX1            : out    vl_logic_vector(6 downto 0);
        HEX2            : out    vl_logic_vector(6 downto 0);
        HEX3            : out    vl_logic_vector(6 downto 0);
        HEX4            : out    vl_logic_vector(6 downto 0);
        HEX5            : out    vl_logic_vector(6 downto 0);
        HEX6            : out    vl_logic_vector(6 downto 0);
        HEX7            : out    vl_logic_vector(6 downto 0);
        State_LED       : out    vl_logic_vector(1 downto 0);
        quick_low_led   : out    vl_logic;
        read_led        : out    vl_logic;
        write_led       : out    vl_logic;
        arload_led      : out    vl_logic;
        arinc_led       : out    vl_logic;
        pcinc_led       : out    vl_logic;
        pcload_led      : out    vl_logic;
        drload_led      : out    vl_logic;
        trload_led      : out    vl_logic;
        irload_led      : out    vl_logic;
        r1load_led      : out    vl_logic;
        r0load_led      : out    vl_logic;
        zload_led       : out    vl_logic;
        pcbus_led       : out    vl_logic;
        drhbus_led      : out    vl_logic;
        drlbus_led      : out    vl_logic;
        trbus_led       : out    vl_logic;
        r1bus_led       : out    vl_logic;
        r0bus_led       : out    vl_logic;
        membus_led      : out    vl_logic;
        busmem_led      : out    vl_logic;
        clr_led         : out    vl_logic
    );
end light_show;
